library ieee;
use ieee.std_logic_1164.all;

package types is
  type mult_arr is array(natural range<>,natural range<>) of std_logic;
end types;
